module led(switch, led);
	input switch;
	output led;
	
	assign led=switch;
endmodule