library verilog;
use verilog.vl_types.all;
entity decorder_tb is
end decorder_tb;
